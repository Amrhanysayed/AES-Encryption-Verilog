module round_inverse(input [127:0]state,input [127:0]key,output wire [127:0]out);
wire[127:0]states[3:0];
InvShiftRows row(state, states[0]);
InvSubBytes SUB(states[0], states[1]);
AddRoundKey k(states[1],key,states[2]);
InvMixColumns inv(states[2],states[3]);
assign out=states[3];

endmodule
module Cipher;

endmodule

module Decipher;

endmodule

module Encrypt  #(parameter nk=4,parameter nr=10) (key);
    input wire [(nk*32)-1:0] key;

endmodule